// maxhpc: Maxim Vorontsov

module ecpix5(
 `include "ecpix5_ports.hv"
);
/* Reset */
 assign rst_sys_ = 1'bz;
/**/

endmodule
